* CMOS Inverter
* BATUHAN TOPALOĞLU 2019 

* SPICE3 file created from nNotEqualt2p.ext - technology: scmos

.option scale=0.12u

*
*TRANSISTOR
*Mname DRAIN GATE SOURCE SUBSTRATE MODEL WIDTH   LENGTH
*      NODE  NODE NODE   NODE      NAME  MICRONS MICRONS
*----- ----- ---- ------ --------- ----  ------- ------
M1000 	y     a   vdd     w_n8_8#  pmos   w=20     l=2
+  ad=100 pd=50 as=100 ps=50

M1001   y     a   gnd      Gnd     nmos   w=8      l=2
+  ad=40 pd=26 as=40 ps=26

*
*CAPACITOR
*Cname +NODE -NODE VALUE(Picofarads)
*----- ----- ----- -----------------
C0 	gnd    y     0.12fF
C1 	gnd    a     0.04fF
C2 	y     vdd    0.25fF
C3	y      a     0.05fF
C4 	y    w_n8_8# 0.07fF
C5 	vdd    a     0.04fF
C6	vdd  w_n8_8# 0.10fF
C7	a    w_n8_8# 0.13fF
C8	gnd   Gnd    0.10fF
C9	y     Gnd    0.05fF
C10	vdd   Gnd    0.02fF
C11	a     Gnd    0.13fF
C12 	w_n8_8# Gnd  0.73fF

*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    vdd    GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     a     GND    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
